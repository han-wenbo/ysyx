import "DPI-C" pure function int  dpi_pmem_read (input int raddr);
import "DPI-C" function void dpi_pmem_write(input int waddr,
                                        input int wdata,
                                        input byte wmask);


module MemContrl(
    input  clk,
    input         valid,
    input         wen,
    input  [31:0] raddr,
    input  [31:0] waddr,
    input  [31:0] wdata,
    input  [7:0]  wmask,
    output reg [31:0] rdata
);

    /* -------- 异步读：组合逻辑 -------- */
    always @(*) begin
        if (valid)
            rdata = dpi_pmem_read(raddr);  // 纯函数，多调无副作用
        else
            rdata = 32'b0;
    end

    /* -------- 同步写：时序逻辑 -------- */
    always @(posedge clk) begin
        if (valid && wen)
            dpi_pmem_write(waddr, wdata, wmask);  // 每拍只执行一次
    end

endmodule
